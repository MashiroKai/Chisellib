module mode (
        input       clk,
        input       rst_n,
        input       mode,
);

endmodule