/*
// 例化 FIFO2Usb_Sync 模块
FIFO2Usb_Sync #(
    .WIDTH(8),                // 设置数据位宽
    .WRFIFO_DEPTH(131072),    // 设置写FIFO深度
    .RDFIFO_DEPTH(512),       // 设置读FIFO深度
    .SENDTHRESHOUD(66048),    // 设置发送阈值
    .WUSEDW(17),              // 设置写使用位宽
    .RUSEDW(9)                // 设置读使用位宽
) my_fifo_usb_sync (
    // 系统接口
    .sys_clk(sys_clk),
    .sys_rst_n(sys_rst_n),
    // FIFO接口
    .VALID(valid_signal),
    .FIFO_DIN(data_in_signal),
    .WR_USEDW(write_used_width_signal),
    .FULL(full_signal),
    .LOAD(load_signal),
    .FIFO_VALID(fifo_valid_signal),
    .FIFO_DOUT(data_out_signal),
    .EMPTY(empty_signal),
    .RD_USEDW(read_used_width_signal),
    // USB模块接口
    .ft232_clk(ft232_clk),
    .ft232_rst_n(ft232_rst_n),
    .D(data_bus),
    .RXF_N(rxf_n_signal),
    .TXE_N(txe_n_signal),
    .RD_N(rd_n_signal),
    .WR_N(wr_n_signal),
    .SIWU_N(siwu_n_signal),
    .OE_N(oe_n_signal)
);

*/


module FIFO2Usb_Sync#(
    // DATA WIDTH AND FIFO DEPTH
    parameter WIDTH = 8,
    parameter WRFIFO_DEPTH = 131072, // WRFIFO DEPTH MUST BIGGER THAN SEND THERSHOLD
    parameter RDFIFO_DEPTH = 512,
    parameter SENDTHRESHOUD = 66048,
    parameter WUSEDW = 17,
    parameter RUSEDW = 9
)
(
    //SYSTEM INTERFACE
     input      sys_clk   
    ,input      sys_rst_n
    //FIFO INTERFACE
    ,input      VALID
    ,input      [WIDTH-1:0]FIFO_DIN
    ,output     [WUSEDW:0]WR_USEDW
    ,output     FULL
    ,input      LOAD        //load data from fifo
    ,output     reg FIFO_VALID     // fifo will output valid and data after 1 clock period if load == 1 and empty == 0; 
    ,output     [WIDTH-1:0]FIFO_DOUT
    ,output     EMPTY
    ,output     [RUSEDW:0]RD_USEDW

    //USB MODULE INTERFACE
    ,input      ft232_clk   //FT232 BOARD 60MHZ CLOCK
    ,input      ft232_rst_n
    ,inout      [WIDTH-1:0]D
    ,input      RXF_N //indicate if the data is avaliable to read from usb fifo
    ,input      TXE_N //indicate if the data can be wirtten to usb fifo 
    ,output     reg RD_N  //usb fifo rd control 
    ,output     reg WR_N  //usb fifo wr control
    ,output     reg SIWU_N  //tie to high
    ,output     reg OE_N  //OUT ENABLE , LOW EFFECTIVE
    // wr/rd one data at a time
);
wire [WIDTH-1:0]DOUT;
assign D= FLAG?DOUT:8'bzzzzzzzz;
// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.


// Generated by Quartus Prime Version 20.1 (Build Build 711 06/05/2020)
// Created on Tue Jan 23 11:29:01 2024

async_fifo_fwft async_fifo_fwft_inst
(
	.data(FIFO_DIN) ,	// input [7:0] data_sig
	.rdclk(ft232_clk) ,	// input  rdclk_sig
	.rdreq(WR_LOAD) ,	// input  rdreq_sig
	.wrclk(sys_clk) ,	// input  wrclk_sig
	.wrreq(VALID) ,	// input  wrreq_sig
	.q(DOUT) ,	// output [7:0] q_sig
	.rdempty(WR_EMPTY) ,	// output  rdempty_sig
	.rdusedw(WR_RD_USEDW) ,	// output [12:0] rdusedw_sig
	.wrfull(FULL) ,	// output  wrfull_sig
	.wrusedw(WR_USEDW) 	// output [12:0] wrusedw_sig
);

reg WR_LOAD;
wire    [logb2(WRFIFO_DEPTH):0]WR_RD_USEDW;
wire    [logb2(WRFIFO_DEPTH):0]RD_WR_USEDW;
async_fifo async_fifo_inst
(
	.data(RD_FIFO_DIN) ,	// input [7:0] data_sig
	.rdclk(sys_clk) ,	// input  rdclk_sig
	.rdreq(LOAD) ,	// input  rdreq_sig
	.wrclk(ft232_clk) ,	// input  wrclk_sig
	.wrreq(RD_FIFO_VALID) ,	// input  wrreq_sig
	.q(FIFO_DOUT) ,	// output [7:0] q_sig
	.rdempty(EMPTY) ,	// output  rdempty_sig
	.rdusedw(RD_USEDW) ,	// output [8:0] rdusedw_sig
	.wrfull(RD_FULL) ,	// output  wrfull_sig
	.wrusedw(RD_WR_USEDW) 	// output [8:0] wrusedw_sig
);
always @(posedge sys_clk or negedge sys_rst_n) begin
    if (!sys_rst_n) begin
        FIFO_VALID <= 1'b0;
    end
    else begin
        FIFO_VALID <= LOAD ;
    end
end
counter #(
    .RST(SENDTHRESHOUD),
    .START(0)
)
sendcnt(
    .clk(ft232_clk)
    ,.rst_n(ft232_rst_n)
    ,.asyn(1'b0)
    ,.en(~WR_N)
    ,.pulse(SEND_CMPLE)
);
wire SEND_CMPLE;
wire RD_FULL;
reg RD_FIFO_VALID;
reg RD_FIFO_DIN;
reg FLAG;
reg [2:0]STATE;
localparam   IDLE = 3'b000;
localparam   RD_STATE_OE_N = 3'b001;
localparam   RD_STATE_RD_N = 3'b010;
localparam   WR_STATE_LOAD = 3'b011;
localparam   WR_STATE_WR_N = 3'b100;
localparam   RD_WAIT = 3'b101;
localparam   WR_WAIT = 3'b110;
always @(posedge ft232_clk or negedge ft232_rst_n) begin
    if (!ft232_rst_n) begin
        STATE <= IDLE;
        FLAG <= 1'b0;
    end
    else begin
        case (STATE)
        IDLE    : begin
                FLAG <= 1'b0;
            if (!RD_FULL&&!RXF_N) begin // RD_FIFO isn't FULL, and there are data avaliable , then read data from FT232
                STATE <= RD_STATE_OE_N;
            end
            else begin
            if (!WR_EMPTY&&!TXE_N&&SEND_ENABLE) begin //WR_FIFO isn't EMPTY,and FT232 is ready to receive data , then write data to FT232
                STATE <= WR_STATE_WR_N;
                FLAG <= 1'b1;
            end
            end
        end
        RD_STATE_OE_N    :begin
                STATE  <=   RD_STATE_RD_N;
        end
        RD_STATE_RD_N    :begin
                if (RD_FULL||RXF_N) begin
                    STATE   <=  IDLE;
                end
        end
        WR_STATE_WR_N    :begin
                if (WR_EMPTY||TXE_N) begin
                    STATE   <=  IDLE;
                end 
        end
        endcase
    end
end
reg SEND_ENABLE;
always @(*) begin
    if (!ft232_rst_n) begin
        SEND_ENABLE <= 1'b0;
    end
    else begin
        if (SEND_CMPLE) begin
            SEND_ENABLE <= 1'b0;
        end
        else begin
            if (WR_RD_USEDW >=SENDTHRESHOUD) begin
            SEND_ENABLE <= 1'b1;
            end
        end
    end
end
always @(*) begin
    if (!ft232_rst_n) begin
        OE_N = 1'b1;
    end
    else begin
        if ((STATE == RD_STATE_OE_N || STATE == RD_STATE_RD_N)&&!RD_FULL&&!RXF_N) begin
            OE_N = 1'b0;
        end
        else begin
            OE_N = 1'b1;
        end
    end
end
always @(*) begin
    if (!ft232_rst_n) begin
        RD_N = 1'b1;
    end
    else begin
        if ((STATE == RD_STATE_RD_N)&&!RD_FULL&&!RXF_N) begin
            RD_N = 1'b0;
        end
        else begin
            RD_N = 1'b1;
        end
    end
end
always @(*) begin
    if (!ft232_rst_n) begin
        WR_N = 1'b1;
    end
    else begin
        if ((STATE == WR_STATE_WR_N )&&!TXE_N&&!WR_EMPTY) begin
            WR_N = 1'b0;
        end
        else begin
            WR_N = 1'b1;
        end
    end
end
always @(*) begin
    if (!ft232_rst_n) begin
        RD_FIFO_VALID = 1'b0;
    end
    else begin
        if ((STATE == RD_STATE_RD_N)&&!RXF_N&&!RD_FULL) begin
            RD_FIFO_VALID = 1'b1;
        end
        else begin
            RD_FIFO_VALID = 1'b0;
        end
    end
end
always @(*) begin
    if (!ft232_rst_n) begin
        WR_LOAD = 1'b0; 
    end
    else begin
        if ((STATE == WR_STATE_WR_N)&&!TXE_N&&!WR_EMPTY) begin
            WR_LOAD = 1'b1;
        end
        else begin
            WR_LOAD = 1'b0;
        end
    end
end

always @(*) begin
    if (!ft232_rst_n) begin
        RD_FIFO_DIN = 8'b0;
    end
    else begin
        if ((STATE == RD_STATE_RD_N)&&!RXF_N&&!RD_FULL) begin
            RD_FIFO_DIN = D;
        end
        else begin
            RD_FIFO_DIN = RD_FIFO_DIN;
        end
    end
end


function integer logb2;
    input [31:0]            value;
    reg   [31:0]            tmp;
begin
    tmp = value - 1;
    for (logb2 = 0; tmp > 0; logb2 = logb2 + 1) 
        tmp = tmp >> 1;
end
endfunction
endmodule
